/* Copyright(C) 2020 Cobac.Net All Rights Reserved. */
/* chapter: ��2��                           */
/* project: blinkspeed                      */
/* outline: LED�̓_�ő��x���v�b�V��SW�Ő��� */

module blinkspeed (
    input               CLK,
    input               RST,
    input       [0:0]   BTN,
    output  reg [2:0]   LED_RGB
);

/* �`���^�����O������H��ڑ� */
wire btnon;

debounce d0 (.CLK(CLK), .RST(RST), .BTNIN(BTN), .BTNOUT(btnon));

/* ���x�ݒ�p�J�E���^ */
reg [1:0] speed;

always @( posedge CLK ) begin
    if ( RST )
        speed <= 2'h0;
    else if ( btnon )
        speed <= speed + 2'h1;
end

/* �V�X�e���N���b�N�𕪎� */
reg [26:0] cnt27;

always @( posedge CLK ) begin
    if ( RST )
        cnt27 <= 27'h0;
    else
        cnt27 <= cnt27 + 27'h1;
end

/* LED�p�J�E���^�̃C�l�[�u�����쐬 */
reg ledcnten;

always @* begin
    case ( speed )
        2'h0:   ledcnten = (cnt27      ==27'h7ffffff);
        2'h1:   ledcnten = (cnt27[25:0]==26'h3ffffff);
        2'h2:   ledcnten = (cnt27[24:0]==25'h1ffffff);
        2'h3:   ledcnten = (cnt27[23:0]==24'hffffff);
        default ledcnten = 1'b0;
    endcase
end

/* LED�p5�i�J�E���^ */
reg [2:0] cnt3;

always @( posedge CLK ) begin
    if ( RST )
        cnt3 <= 3'h0;
    else if ( ledcnten )
        if ( cnt3==3'd4)
            cnt3 <=3'h0;
        else
            cnt3 <= cnt3 + 3'h1;
end

/* LED�f�R�[�_ */
always @* begin
    case ( cnt3 )
        3'd0:   LED_RGB = 3'b100;
        3'd1:   LED_RGB = 3'b010;
        3'd2:   LED_RGB = 3'b001;
        3'd3:   LED_RGB = 3'b111;
        3'd4:   LED_RGB = 3'b000;
        default:LED_RGB = 3'b000;
    endcase
end

endmodule